`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/12/15 16:37:49
// Design Name: 
// Module Name: simple_column_scanner_pipeline
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module simple_column_scanner_pipeline #(
  parameter integer OUT_W   = 112,
  parameter integer OUT_H   = 112,
  parameter integer TILE_H  = 6,
  parameter integer COUT    = 32,
  parameter integer UNIT_NUM= 16,
  parameter integer K       = 3,
  parameter integer PADDING = 1
)(
  input  wire clk,
  input  wire rst_n,

  // ���������źţ�ÿ�� batch ������һ�ļ���
  input  wire start,

  // Prefetch ����
  output reg  prefetch_start,
  output reg  [$clog2(OUT_H)-1:0] prefetch_tile_row,
  input  wire prefetch_done,
  input  wire prefetch_busy,
  input  wire buffer_ready,

  // ��������
  output wire read_enable,
  output wire [$clog2(OUT_W+2*PADDING)-1:0] read_addr,

  // ״ָ̬ʾ
  output reg  busy,
  output reg  done,
  output reg  [$clog2(OUT_W+2*PADDING)-1:0] current_col
);

  // ���β���
  localparam integer STRIDE    = TILE_H - K + 1;
  localparam integer PADDED_W  = OUT_W + 2 * PADDING;
  localparam integer PADDED_H  = OUT_H + 2 * PADDING;
  localparam integer NUM_TILES = (PADDED_H - TILE_H) / STRIDE + 1;

  // ״̬��
  localparam IDLE          = 3'd0;
  localparam PREFETCH_FIRST= 3'd1;
  localparam SCAN          = 3'd2;
  localparam DONE_ST       = 3'd3;

  reg [2:0] state;

  reg [$clog2(NUM_TILES)-1:0] scan_tile_idx;
  reg [$clog2(PADDED_W)-1:0]  col_counter;

  // FSM
  always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      state            <= IDLE;
      scan_tile_idx    <= 0;
      col_counter      <= 0;
      prefetch_start   <= 0;
      prefetch_tile_row<= 0;
      busy             <= 0;
      done             <= 0;
      current_col      <= 0;
    end else begin
      // Ĭ��������
      prefetch_start <= 0;
      done           <= 0;

      // start ��Ϊ�����ȼ���λ�����۵�ǰ��ʲô״̬����һ�� start �ʹ�ͷ��ʼɨ��
      if (start) begin
        busy             <= 1'b1;
        state            <= PREFETCH_FIRST;
        scan_tile_idx    <= 0;
        col_counter      <= 0;
        prefetch_tile_row<= 0;
        prefetch_start   <= 1'b1;   // ������һ�� tile ��Ԥȡ
      end else begin
        case (state)
          IDLE: begin
            busy <= 1'b0;
            // ��������ȴ� start����Ϊ�����Ѿ������� start ��֧
          end

          PREFETCH_FIRST: begin
            // �ȴ� prefetch_double_buffer �ѵ�ǰ tile ����
            if (prefetch_done && buffer_ready) begin
              col_counter <= 0;
              state       <= SCAN;
            end
          end

          SCAN: begin
            // һ��һ�е�ɨ�赱ǰ tile
            current_col <= col_counter;

            if (col_counter < PADDED_W-1) begin
              col_counter <= col_counter + 1'b1;
            end else begin
              // ��ǰ tile ��һ��ɨ�����
              if (scan_tile_idx < NUM_TILES-1) begin
                // ������һ tile ��
                scan_tile_idx    <= scan_tile_idx + 1'b1;
                col_counter      <= 0;
                prefetch_tile_row<= prefetch_tile_row + STRIDE;
                prefetch_start   <= 1'b1;
                state            <= PREFETCH_FIRST;
              end else begin
                // ���� tile ɨ�����
                state <= DONE_ST;
              end
            end
          end

          DONE_ST: begin
            busy <= 1'b0;
            done <= 1'b1;   // �� done һ��
            state <= IDLE;
          end

          default: begin
            state <= IDLE;
          end
        endcase
      end
    end
  end

  // ��ʹ�� / ��ַ��ֻҪ�� SCAN ״̬���� buffer_ready���Ϳ��Դ� prefetch buffer ����Ӧ��
  assign read_enable = (state == SCAN) && buffer_ready;
  assign read_addr   = col_counter;

endmodule