`ifndef MOBILENET_DEFINES_VH
`define MOBILENET_DEFINES_VH

// ============================================================
// MobileNetV1 ȫ�ֲ�������
// ============================================================

// ����λ��
`define DATA_W          8
`define ACC_W           32
`define PSUM_W          18
`define PROD_W          16

// PE��������
`define NUM_ROWS        16
`define NUM_COLS        16
`define UNIT_NUM        16
`define LANES           16

// MobileNetV1 ��������
`define TOTAL_LAYERS    28
`define TOTAL_CONV_DW_PW_LAYERS 27  // ����FC

// ���ߴ�����
`define MAX_IMG_W       224
`define MAX_IMG_H       224
`define MAX_CHANNELS    1024
`define MAX_OUT_W       112
`define MAX_OUT_H       112

// ����ͼ�������� (112*112*64 / 16 = 50176 words)
`define FEATURE_BUF_DEPTH   50176

// Ȩ�ش洢����ַ (Layer0��0��ʼ, Layer2��64��ʼ)
`define L0_WEIGHT_BASE      9'd0
`define L2_WEIGHT_BASE      9'd64

// ����·�� (����ʵ�ʻ����޸�)
`define DATA_PATH           "D:/NoC/mycode/mobilenet_acc2/data/"

// ============ Layer Type Definitions (3-bit) ============
localparam [2:0] LAYER_TYPE_CONV = 3'd0;  // ��һ���׼3x3���
localparam [2:0] LAYER_TYPE_DW   = 3'd1;  // Depthwise Convolution
localparam [2:0] LAYER_TYPE_PW   = 3'd2;  // Pointwise Convolution
localparam [2:0] LAYER_TYPE_AP   = 3'd3;  // Global Average Pooling
localparam [2:0] LAYER_TYPE_FC   = 3'd4;  // Fully Connected

// ============ MobileNetV1 Layer Count ============
localparam integer TOTAL_LAYERS = 29;  // Layer 0-28 (��29��)
localparam integer MAX_LAYER_ID = 28;  // ���һ��ID

// ============ Data Width ============
localparam integer DATA_W    = 8;      // INT8
localparam integer ACC_W     = 32;     // �ۼ���λ��
localparam integer WEIGHT_W  = 8;      // Ȩ��λ��

// ============ PE Array Size ============
localparam integer PE_ROWS   = 16;
localparam integer PE_COLS   = 16;

// ============ Memory Parameters ============
localparam integer WEIGHT_ADDR_W = 16;
localparam integer BIAS_ADDR_W   = 12;
localparam integer FEAT_ADDR_W   = 17;

`endif